
------------------------------------------------------------------------
-- VGA Display demo code
-- Numato Lab
-- http://www.numato.com
-- http://www.numato.cc
-- License : CC BY-SA (http:-creativecommons.org/licenses/by-sa/2.0/)
-------------------------------------------------------------------------

library IEEE;
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity VGADisplay is
    -- Define the width and the height of the displayed text.
		generic(OutputWidth: integer := 10;	  
			   OutputHeight: integer := 40	 
			   );
		  port (
	-- Assuming 50MHz clock.If the clock is reduced then it might give the unexpected output.	   
			  clock: in std_logic;
			  Switch: in std_logic_vector(5 downto 0);
			  
	-- The counter tells whether the correct position on the screen is reached where the data is to be displayed. 
			  hcounter: in integer range 0 to 1023;
			  vcounter: in integer range 0 to 1023;
	
	-- Output the colour that should appear on the screen. 
			  pixels : out std_logic_vector(7 downto 0)				  
			  );
end VGADisplay;


architecture Behavioral of VGADisplay is	
    -- Intermediate register telling the exact position on display on screen.
		 signal game_over : std_logic := '0';
		 signal explosion : integer range 0 to 7 := 0;
		 
		 signal x : integer range 0 to 640 := 640;
		 signal y : integer range 0 to 480 := 124;
		 signal row : std_logic_vector(47 downto 0);
		 
		 
		 signal x2 : integer range 0 to 640 := 640;
		 signal y2 : integer range 0 to 480 := 224;
		 signal row2 : std_logic_vector(47 downto 0);
		 
		 signal x3 : integer range 0 to 640 := 640;
		 signal y3 : integer range 0 to 480 := 324;
		 signal row3 : std_logic_vector(47 downto 0);
		 
		 signal xS : integer range 0 to 640 := 30;
		 signal yS : integer range 0 to 480 := 224;
		 signal rowS : std_logic_vector(47 downto 0);
		 
		 signal xG : integer range 0 to 640 := 296;
		 signal yG : integer range 0 to 480 := 216;
		 signal rowG : std_logic_vector(47 downto 0);
		 
		 signal animate_counter_x : std_logic_vector(30 downto 0) := (others => '0');
		 signal animate_counter_y : std_logic_vector(30 downto 0) := (others => '0');
		 
		 signal debounce_counter_up : integer range 0 to 5 := 0;
		 signal debounce_counter_down : integer range 0 to 5 := 0;

		 signal meteor_spawn_delay_counter : integer range 0 to 300 := 0;
		 signal spawn_meteor1 : std_logic := '0';
		 signal spawn_meteor2 : std_logic := '0';
		 signal spawn_meteor3 : std_logic := '0';
		 
		 signal ship_anim_counter : integer range 0 to 3 := 0;
		 
	type font is array (0 to 47) of std_logic_vector(47 downto 0);

signal game_over_graphic : font := (
"000000000000000000000000000000000000000000000000",
"000000000000000000000000000000000000000000000000",
"000000000000000000000000000000000000000000000000",
"000000000000000000000000000000000000000000000000",
"000000000000000000000000000000000000000000000000",
"000000000000000000000000000000000000000000000000",
"000000000000000000000000000000000000000000000000",
"000000000000000000000000000000000000000000000000",
"000000000000000000000000000000000000000000000000",
"000000000000000000000000000000000000000000000000",
"000000000000000000000000000000000000000000000000",
"000000000000000000000000000000000000000000000000",
"000000000000000000000000000000000000000000000000",
"000000000000000000000000000000000000000000000000",
"000000111111100110000110000111000011111100000000",
"000000000001100111001110001101100000000110000000",
"000000000001100111111110011000110000000011000000",
"000000000001100111111110111000111000000011100000",
"000000111111100110100110111000111011110011100000",
"000000000001100110000110111111111011000011100000",
"000000000001100110000110111000111011000110000000",
"000000111111100110000110111000111011111100000000",
"000000111111100110000110010000010011111100000000",
"000000000000000000000000000000000000000000000000",
"000000011111111011111110111000111001111110000000",
"000000110000111000000110111000111011100011000000",
"000000110000111000000110111000111011000011100000",
"000000111000111000001110111000111011000011100000",
"000000111100111011111110111101111011000011100000",
"000000001111111000000110001111110011000011100000",
"000000011110111000000110000111000011000011100000",
"000000111100111011111110000010000001111111000000",
"000000000000000000000000000000000000000000000000",
"000000000000000000000000000000000000000000000000",
"000000000000000000000000000000000000000000000000",
"000000000000000000000000000000000000000000000000",
"000000000000000000000000000000000000000000000000",
"000000000000000000000000000000000000000000000000",
"000000000000000000000000000000000000000000000000",
"000000000000000000000000000000000000000000000000",
"000000000000000000000000000000000000000000000000",
"000000000000000000000000000000000000000000000000",
"000000000000000000000000000000000000000000000000",
"000000000000000000000000000000000000000000000000",
"000000000000000000000000000000000000000000000000",
"000000000000000000000000000000000000000000000000",
"000000000000000000000000000000000000000000000000",
"000000000000000000000000000000000000000000000000"
);

signal m : font := (
"000000000000000000000000000000000000000000000000",
"000000000000000000000011100000000000000000000000",
"000000000000000011111100110000000000000000000000",
"000000000000001111110000001100000000000000000000",
"000000000000111110000000000100000000000000000000",
"000000000011111100000000000010000000000000000000",
"000000011111111100000000000011000000000000000000",
"000001111111111111000000000011111000000000000000",
"000011111111111111110000000011111110000000000000",
"000111111111111111111000011100011111110000000000",
"001111111111111111111000110000000000111100000000",
"011111111111111111111100110000000000000111100000",
"011111111111111111111111110000000000000001100000",
"011111111111111111111111110000000000000000110000",
"011111111101111111111111110000000000000000110000",
"011111111110000001111111111000000000000000110000",
"011111111111000001111111111000000000000000010000",
"011111111111111000111111111100011000000000010000",
"011111111111111000111111111111111110000000111000",
"011111111111111111111111111111111111000011111000",
"011111111111111111111111111111111111000011111000",
"011111111111111111111111111111111110000000011000",
"001111111111111111111111111111111110000000001000",
"001111111111111111111111111111111110000000001100",
"001111111111111111111111111111111111000000000100",
"001111111111111111111111111111111111111111000010",
"001111111111111111111111111111110011111111100000",
"000111111111111111111111111111110000000011111010",
"000011111111111111111111111111110000000000011110",
"000000111111111111111111111111110000000000011110",
"000000011111111111111111111111111000000000011110",
"000000001111111111111111111111111100000000011100",
"000000000011111111111111111001111100000000111000",
"000000000001111111111111111001111110000011110000",
"000000000000001111111111111101111111111111000000",
"000000000000000111111111111101111111111110000000",
"000000000000000111111111111100111111111100000000",
"000000000000000011111111111111111111111100000000",
"000000000000000011111111111111111111111100000000",
"000000000000000011111111111111111111111000000000",
"000000000000000001111111111111111111111000000000",
"000000000000000001111111111111111111111000000000",
"000000000000000000011111111111111111111000000000",
"000000000000000000000001111111111111111000000000",
"000000000000000000000000001111111111110000000000",
"000000000000000000000000000001111111110000000000",
"000000000000000000000000000000000000000000000000",
"000000000000000000000000000000000000000000000000"
);
		
signal m2 : font := (
"000000000000000000000000000000000000000000000000",
"000000000000000000000000000000000000000000000000",
"000000000000000000000000000000000000000000000000",
"000000000000000000000000000000011100000000000000",
"000000000000000000000001111111100100000000000000",
"000000000000000111111111000000000010000000000000",
"000000000000111111111110000000000011000000000000",
"000000000001100000000000000000000001000000000000",
"000000000111000000000000000000000000100000000000",
"000000011100000000000000000000000000110000000000",
"000000111000000000000000010000000000010000000000",
"000000111100000111000000010000000000011000000000",
"000000111111111111111000010000000000001000000000",
"000000111111111111111111110000000000001100000000",
"000001111111111101111111110000000000100110000000",
"000001011111111100111111110000000000111111000000",
"000011001111111100011111110000000000111111000000",
"000011000111111100001111110000000000111001100000",
"000111000111111110000001111000000000111100010000",
"000111111111111111100011111100000000011110001000",
"000111111111111111111110001100000000001111001000",
"001111111111111111111000000110000000001111001000",
"000111111111111111111111110011000000000111001000",
"000111111111111111111111111111111111111111001100",
"000111111111111111111111111111111111111111100100",
"001111111111111111111111111111111111111111110100",
"001111111111111111111111111111111111111111111000",
"001111111111111111111111111111111111111111111110",
"011111111111111111111111111111111111110011111110",
"011111111111111111011111111111111111100011111110",
"001111111111111111000000111111111111000011111100",
"000111111111111111000000011111111111000000111100",
"000111111111111111000000001111111111111110011000",
"000011111111111111110000000000111111111111111000",
"000001111111111111111100000111111111111111110000",
"000001111111111111111111111111111111111111110000",
"000000111111111111111111111111111111111111110000",
"000000011111111111111111111111111111111111100000",
"000000001111111111111111111111111111111111100000",
"000000001111111111111111111111111111111111000000",
"000000000111111111111111111111111111111111000000",
"000000000011111101111111111111111100000000000000",
"000000000001000000000111111111100000000000000000",
"000000000000000000000000011100000000000000000000",
"000000000000000000000000000000000000000000000000",
"000000000000000000000000000000000000000000000000",
"000000000000000000000000000000000000000000000000",
"000000000000000000000000000000000000000000000000"
);

signal m3 : font := (
"000000000000000000000000000000000000000000000000",
"000000001000000000000000000000000000000000000000",
"000000011111100000110000000000000000000000000000",
"000000111111111111111100000000000000000000000000",
"000001111111111111111110000000000000000000000000",
"000011111111111111110001000000000000000000000000",
"000111111111111111111000000000000000000000000000",
"001111111111111111101111111100000000000000000000",
"011111111111111111000111111000000000000000000000",
"011111111111111111001111111000000000000000000000",
"001111111111111111101111111000000000000000000000",
"000111111111111111100111111000000000000000000000",
"000111111111111111000111111000000000000000000000",
"000011111111111111001111000000000010000000000000",
"000011111111111111001110000000000010000000000000",
"000011111111111111011110000000000011000000000000",
"000011111111111111111110000000000011000000000000",
"000011111111111111111110000000000011000000000000",
"000011111111111111111100000000000011100000000000",
"000011111111111111111100000000000010111000000000",
"000011111111111111111100000000000010000110000000",
"000011111111111111111100000000000111000011100000",
"000011111111111111100000000001111111000001010000",
"000011111111111111100000000011111111000000001000",
"000011111111111111100000000111111111000000000100",
"000011111111111111000000000110000111000000000100",
"000011111111111111100000011110000000000000000000",
"000011111111111111100111111100000000000000000000",
"000011111111111111111111111100000000000000000000",
"000011111111111111111111111000000000110000000000",
"000001111111111111111111111000000001100000000000",
"000001111111111111111111111100000001000000000000",
"000000111111111111111111111110000111000000000000",
"000000111111111111111111111111001111000000000000",
"000000011111111111111111111111111111100000000000",
"000000001111111111111111111111111111100000000000",
"000000000111111111111111111111111111110000000000",
"000000000011111111111111111111111111110010000000",
"000000000001111111111111111111111111111111100100",
"000000000000111000111111111111111110001111111100",
"000000000000000000011111111111111100001111000000",
"000000000000000000000111111111111110001110000000",
"000000000000000000000011111111111110001000000000",
"000000000000000000000000111111111110000000000000",
"000000000000000000000000011111111110000000000000",
"000000000000000000000000000001111110000000000000",
"000000000000000000000000000000001100000000000000",
"000000000000000000000000000000000000000000000000"
);

signal ho229_flight_unit1 : font := (
"000000000000000000000000000000000000000000000000",
"000000000000011000000000000000000000000000000000",
"000000000001110000000000000000000000000000000000",
"000000000000110000000000000000000000000000000000",
"000000000000011000000000000000000000000000000000",
"000000000000001110000000000000000000000000000000",
"000000000000001111000000000000000000000000000000",
"000000000000000111100000000000000000000000000000",
"000000000000000011111000000110000000000000000000",
"000000000000000001111100001100000000000000000000",
"000000000000011111111110011100000000000000000000",
"000000000000111111111111111100000000000000000000",
"000000000000111111111111011100000000000000000000",
"000000000000001111111111000000000000000000000000",
"000000000000000111110000000000000000000000000000",
"000000000000000111100000000000000000000000000000",
"000000000000001111100010000000000000000000000000",
"000000000000011111100110000000000000000000000000",
"000000000000111111001110000000000000000000000000",
"000000000001111111111111111100100000000000000000",
"000000000011001111111111111100100000000000000000",
"000000000111001111111110000000000000000000000000",
"000000001111001111111111110000000000000000000000",
"000000111111111111111111111111111111111100000000",
"000000111111111111111111111111111111111100000000",
"000000001111001111111111110000000000000000000000",
"000000000111001111111110000000000000000000000000",
"000000000011001111111111111100100000000000000000",
"000000000001111111111111111100100000000000000000",
"000000000000111111001110000000000000000000000000",
"000000000000011111100110000000000000000000000000",
"000000000000001111100010000000000000000000000000",
"000000000000001111100000000000000000000000000000",
"000000000000000111110000000000000000000000000000",
"000000000000001111111111000000000000000000000000",
"000000000000111111111111011100000000000000000000",
"000000000000111111111111111100000000000000000000",
"000000000000011111111110011100000000000000000000",
"000000000000000001111100001100000000000000000000",
"000000000000000011111000000110000000000000000000",
"000000000000000111100000000000000000000000000000",
"000000000000001111000000000000000000000000000000",
"000000000000001110000000000000000000000000000000",
"000000000000011000000000000000000000000000000000",
"000000000000110000000000000000000000000000000000",
"000000000001110000000000000000000000000000000000",
"000000000000011000000000000000000000000000000000",
"000000000000000000000000000000000000000000000000"
);
signal ho229_flight_unit2 : font := (
"000000000000000000000000000000000000000000000000",
"000000000000011000000000000000000000000000000000",
"000000000001110000000000000000000000000000000000",
"000000000000110000000000000000000000000000000000",
"000000000000011000000000000000000000000000000000",
"000000000000001110000000000000000000000000000000",
"000000000000001111000000000000000000000000000000",
"000000000000000111100000000000000000000000000000",
"000000000000000011111000000110000000000000000000",
"000000000000000001111100001100000000000000000000",
"000000000000011111111110011100000000000000000000",
"000000000000111111111111111100000000000000000000",
"000000000000111111111111011100000000000000000000",
"000000000000001111111111000000000000000000000000",
"000000000000000111110000000000000000000000000000",
"000000000000000111100000000000000000000000000000",
"000000000000001111100010000000000000000000000000",
"000000000000011111100110000000000000000000000000",
"000000000000111111001110000000000111110000000000",
"000000000001111111111111111100101111111111100000",
"000000000011001111111111111100101111111111100000",
"000000000111001111111110000000000111110000000000",
"000000001111001111111111110000000000000000000000",
"000000111111111111111111111111111111111100000000",
"000000111111111111111111111111111111111100000000",
"000000001111001111111111110000000000000000000000",
"000000000111001111111110000000000111110000000000",
"000000000011001111111111111100101111111111100000",
"000000000001111111111111111100101111111111100000",
"000000000000111111001110000000000111110000000000",
"000000000000011111100110000000000000000000000000",
"000000000000001111100010000000000000000000000000",
"000000000000001111100000000000000000000000000000",
"000000000000000111110000000000000000000000000000",
"000000000000001111111111000000000000000000000000",
"000000000000111111111111011100000000000000000000",
"000000000000111111111111111100000000000000000000",
"000000000000011111111110011100000000000000000000",
"000000000000000001111100001100000000000000000000",
"000000000000000011111000000110000000000000000000",
"000000000000000111100000000000000000000000000000",
"000000000000001111000000000000000000000000000000",
"000000000000001110000000000000000000000000000000",
"000000000000011000000000000000000000000000000000",
"000000000000110000000000000000000000000000000000",
"000000000001110000000000000000000000000000000000",
"000000000000011000000000000000000000000000000000",
"000000000000000000000000000000000000000000000000"
);

signal xwing_star_fighter : font := (
"000000000000000000000000000000000000000000000000",
"000000000000000000000000000000000000000000000000",
"000000000000000000000000000000000000000000000000",
"000000000000000000000000000000000000000000000000",
"000000000000000000000000000000000111111000000000",
"000000000000000000000111111111111111111100000000",
"000000000000000000000111111111111111111100000000",
"000000000000000000000000000000000111111000000000",
"000000000000000000000000000000000111111000000000",
"000000000000000000000000000000000111111000000000",
"000000000000000000000000000000000111111000000000",
"000000000000000000000000000000000111111100000000",
"000000000000000000000000000000000111111100000000",
"000000000000000000000000000000000111111100000000",
"000000000000000000000000000000000111111110000000",
"000000000000000000000000000000000111111110000000",
"000000000000000000000000000000000111111110000000",
"000000000000000000000000000000001111111110000000",
"000000000000000000000000000000011111111111111100",
"000000000000000000000000000000011111111111111100",
"000000000000000000000000000000001111111110000000",
"000000000000000000000000000000111111111111000000",
"000000000000000011111111111111111111111111100000",
"001111111111111111110000011111000111111111100000",
"111100111111111110000000001110000011111111100000",
"001111111111111111110000011111000111111111100000",
"000000000000000111111111111111111111111111100000",
"000000000000000000000000000000111111111111000000",
"000000000000000000000000000000001111111110000000",
"000000000000000000000000000000011111111111111100",
"000000000000000000000000000000011111111111111100",
"000000000000000000000000000000001111111110000000",
"000000000000000000000000000000000111111110000000",
"000000000000000000000000000000000111111110000000",
"000000000000000000000000000000000111111110000000",
"000000000000000000000000000000000111111100000000",
"000000000000000000000000000000000111111100000000",
"000000000000000000000000000000000111111100000000",
"000000000000000000000000000000000111111000000000",
"000000000000000000000000000000000111111000000000",
"000000000000000000000000000000000111111000000000",
"000000000000000000000000000000000111111000000000",
"000000000000000000000111111111111111111100000000",
"000000000000000000000111111111111111111100000000",
"000000000000000000000000000000000111111000000000",
"000000000000000000000000000000000000000000000000",
"000000000000000000000000000000000000000000000000",
"000000000000000000000000000000000000000000000000"
);

begin

 -- On every positive edge of the clock counter condition is checked,
  output1: process(clock)
			  begin
			  if rising_edge (clock) then
			  
			  -- Reset Logic
					if (switch(0) = '0') then
						explosion <= 0;
						game_over <= '0';
						x <= 640;
						x2 <= 640;
						x3 <= 640;
						yS <= 224;
						animate_counter_x <= (others => '0');
						animate_counter_y <= (others => '0');
						meteor_spawn_delay_counter <= 0;
						spawn_meteor1 <= '0';
						spawn_meteor2 <= '0';
						spawn_meteor3 <= '0';
					end if;
			  
				 animate_counter_x <= std_logic_vector(unsigned(animate_counter_x) + 1);
				 animate_counter_y <= std_logic_vector(unsigned(animate_counter_y) + 1);
				 if explosion < 7 then
					 if animate_counter_x(20) = '1' then
						
						-- Ship Animation

						ship_anim_counter <= ship_anim_counter + 1;
						
						-- Explosion Timer
						if game_over = '1' and explosion < 7 then
							explosion <= explosion + 1;
						end if;

						-- Meteor Movement
						case spawn_meteor1 is
							when '1' =>
								x <= x - 5;
							when others =>
						end case;
						case spawn_meteor2 is
							when '1' =>
								x2 <= x2 - 3;
							when others =>
						end case;
						case spawn_meteor3 is
							when '1' =>
								x3 <= x3 - 4;
							when others =>
						end case;
--						if spawn_meteor1 = '1' then                      -- replaced with case
--							x <= x - 5;
--						end if ;
--
--						if spawn_meteor2 = '1' then
--							x2 <= x2 - 3;
--						end if ;
--
--						 if spawn_meteor3 = '1' then
--							x3 <= x3 - 4;
--						 end if ;

						-- Delaying the spawns of meteors
						 meteor_spawn_delay_counter <= meteor_spawn_delay_counter + 1;
						 case meteor_spawn_delay_counter is
						 	when 300 => spawn_meteor3 <= '1';
							when 260 => spawn_meteor1 <= '1';
							when 230 => spawn_meteor2 <= '1';
							when others =>
						 end case;
--						 if meteor_spawn_delay_counter = 300 then          --replaced with case
--								spawn_meteor3 <= '1';
--							elsif meteor_spawn_delay_counter = 260 then
--								spawn_meteor1 <= '1';
--							elsif meteor_spawn_delay_counter = 230 then
--								spawn_meteor2 <= '1';
--						 end if ;
						 
						 --Press Switch(2) to move the ship up
						 if (Switch(2) = '0' and yS > 124) then
								debounce_counter_up <= debounce_counter_up + 1;
								case debounce_counter_up is
									when 1 => yS <= yS - 100;
									when others =>
								end case;
								--if debounce_counter_up = 1 then         -- replaced with case
								--	yS <= yS - 100;
								--end if;
						 else
							debounce_counter_up <= 0;
						 end if;
						 
						 --Press Switch(4) to move the ship down
						 if (Switch(4) = '0' and yS < 324) then
								debounce_counter_down <= debounce_counter_down + 1;
								case debounce_counter_down is
									when 1 => yS <= yS + 100;
									when others =>
								end case;
								--if debounce_counter_down = 1 then        -- replaced with case
								--	yS <= yS + 100;
								--end if;
						 else
							debounce_counter_down <= 0;
						 end if;
						 
						 animate_counter_x <= (others => '0');
					 end if;
					 
						-- Meteor vertical movement, Unused
					 if animate_counter_y(20) = '1' then
						 y <= y + 0;
						 y2 <= y2 + 0;
						 y3 <= y3 + 0;
						 animate_counter_y <= (others => '0');
					 end if;

						-- If the counter satisfy the condition, then output the colour that should appear.

						
						-- Checking to see if current pixel is in the ship
						if ship_anim_counter > 2 then
								rowS <= ho229_flight_unit1(vcounter - yS);																		-- SHIP ANIMATION
						else
								rowS <= ho229_flight_unit2(vcounter - yS);
						end if;
						if  (hcounter >= xS and hcounter <= xS + 47 and vcounter >= yS and vcounter <= yS + 47 and rowS(hcounter - xS) = '1') then
								pixels <= x"DB";
							  
						-- Checking to see if current pixel is in object 1
					   elsif  (hcounter >= x and hcounter <= x + 47 and vcounter >= y and vcounter <= y + 47) then
							  row <= m(vcounter - y);
							  if (row(hcounter - x) = '1') then
									pixels <= x"92";
							  else
									pixels <= x"00";
							  end if;
						
						-- Checking to see if current pixel is in object 2
						elsif  (hcounter >= x2 and hcounter <= x2 + 47 and vcounter >= y2 and vcounter <= y2 + 47) then
							  row2 <= m2(vcounter - y2);
							  if (row2(hcounter - x2) = '1') then
									pixels <= x"B7";
							  else
									pixels <= x"00";
							  end if;
						
						-- Checking to see if current pixel is in object 3
						elsif  (hcounter >= x3 and hcounter <= x3 + 47 and vcounter >= y3 and vcounter <= y3 + 47) then
							  row3 <= m3(vcounter - y3);
							  if (row3(hcounter - x3) = '1') then
									pixels <= x"BE";
							  else
									pixels <= x"00";
							  end if;
						
						-- If the condition is not satisfied then the output colour will be black.
						else
							pixels <= x"00";
						end if;
						
						-- Collision Logic
						if yS = y and x >= 47 and x <= 77 then
								game_over <= '1';
						elsif yS = y2 and x2 >= 47 and x2 <= 77 then
								game_over <= '1';
						elsif yS = y3 and  x3 >= 47 and x3 <= 77 then
								game_over <= '1';
						end if;
						
						
						-- Game over screen
					elsif explosion = 7 then
							if  (hcounter >= xG and hcounter <= xG + 47 and vcounter >= yG and vcounter <= yG + 47) then
							  rowG <= game_over_graphic(vcounter - yG);
							  if (rowG(hcounter - xG) = '1') then
									pixels <= x"E0";
							  else
									pixels <= x"00";
							  end if;
							else
								pixels <= x"00";
							end if;
					end if;
			  end if;
		   end process;
			
end Behavioral;
